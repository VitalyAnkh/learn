conectix             $�}vbox   Wi2k     �       �  -   ����A}!
x�@��0s_�0                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������                 ���r                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            conectix             $�}vbox   Wi2k     �       �  -   ����A}!
x�@��0s_�0                                                                                                                                                                                                                                                                                                                                                                                                                                            